module pow_5_pipe_struct
# (
    parameter w = 8
)
(
    input                clk,
    input                rst_n,
    input                n_vld,
    input  [w     - 1:0] n,
    output [        3:0] res_vld,
    output [w * 4 - 1:0] res
);

    wire           n_vld_q_1;
    wire [w - 1:0] n_q_1;

    reg_rst_n        i0_n_vld   (clk, rst_n, n_vld, n_vld_q_1);
    reg_no_rst # (w) i0_n       (clk, n, n_q_1);

    //------------------------------------------------------------------------

    wire [w - 1:0] mul_d_1 = n_q_1 * n_q_1;

    wire           n_vld_q_2;
    wire [w - 1:0] n_q_2;
    wire [w - 1:0] mul_q_2;

    reg_rst_n        i1_n_vld ( clk , rst_n  , n_vld_q_1 , n_vld_q_2 );
    reg_no_rst # (w) i1_n     ( clk ,          n_q_1     , n_q_2     );
    reg_no_rst # (w) i1_mul   ( clk ,          mul_d_1   , mul_q_2   );

    assign res_vld [3]   = n_vld_q_2;
    assign res     [31:24] = mul_q_2;
    
    //------------------------------------------------------------------------

    wire [w - 1:0] mul_d_2 = mul_q_2 * n_q_2;

    wire           n_vld_q_3;
    wire [w - 1:0] n_q_3;
    wire [w - 1:0] mul_q_3;

    reg_rst_n        i2_n_vld ( clk , rst_n  , n_vld_q_2 , n_vld_q_3 );
    reg_no_rst # (w) i2_n     ( clk ,          n_q_2     , n_q_3     );
    reg_no_rst # (w) i2_mul   ( clk ,          mul_d_2   , mul_q_3   );

    assign res_vld [2]     = n_vld_q_3;
    assign res     [23:16] = mul_q_3;

    //------------------------------------------------------------------------

    wire [w - 1:0] mul_d_3 = mul_q_3 * n_q_3;

    wire           n_vld_q_4;
    wire [w - 1:0] n_q_4;
    wire [w - 1:0] mul_q_4;

    reg_rst_n        i3_n_vld ( clk , rst_n  , n_vld_q_3 , n_vld_q_4 );
    reg_no_rst # (w) i3_n     ( clk ,          n_q_3     , n_q_4     );
    reg_no_rst # (w) i3_mul   ( clk ,          mul_d_3   , mul_q_4   );

    assign res_vld [1]    = n_vld_q_4;
    assign res     [15:8] = mul_q_4;

    //------------------------------------------------------------------------

    wire [w - 1:0] mul_d_4 = mul_q_4 * n_q_4;

    wire           n_vld_q_5;
    wire [w - 1:0] n_q_5;
    wire [w - 1:0] mul_q_5;

    reg_rst_n        i4_n_vld ( clk , rst_n  , n_vld_q_4 , n_vld_q_5 );
    reg_no_rst # (w) i4_n     ( clk ,          n_q_4     , n_q_5     );
    reg_no_rst # (w) i4_mul   ( clk ,          mul_d_4   , mul_q_5   );

    assign res_vld [0]   = n_vld_q_5;
    assign res     [7:0] = mul_q_5;

endmodule
