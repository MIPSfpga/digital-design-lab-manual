module pow_5_multi_cycle_always
# (
    parameter w = 8
)
(
    input            clk,
    input            rst_n,
    input            n_vld,
    input  [w - 1:0] n,
    output           res_vld,
    output [w - 1:0] res
);

    reg           n_vld_q;
    reg [w - 1:0] n_q;

    always @ (posedge clk or negedge rst_n)
        if (! rst_n)
            n_vld_q <= 1'b0;
        else
            n_vld_q <= n_vld;

    always @ (posedge clk)
        n_q <= n;

    reg [4:0] shift;

    always @ (posedge clk or negedge rst_n)
        if (! rst_n)
            shift <= 5'b0;
        else if (n_vld_q)
            shift <= 5'b10000;
        else
            shift <= shift >> 1;

    assign res_vld = shift [0];

    reg [w - 1:0] mul;

    always @(posedge clk)
        if (n_vld_q)
            mul <= n_q;
        else
            mul <= mul * n_q;

    assign res = mul;

endmodule
